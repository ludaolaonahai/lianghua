module top;
initial begin
$get_hier();
end
endmodule
