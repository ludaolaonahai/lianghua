module top;
function void myfunc ();
//void'($display(""));
endfunction
endmodule
